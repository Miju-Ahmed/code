module b2e3(e,b);
input[3:0]b;
output[3:0]e;

not(e[0],b[0]);

xnor(e[1],b[1],b[0]);

wire a,c;
or(a,b[0],b[1]);
xor(e[2],b[2],a);

and(c,b[2],a);
or(e[3],b[3],c);
endmodule

