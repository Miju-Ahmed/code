module rc2(j,k,clk,clr,q,qbar);
input j,k,clk,clr;
output[3:0]q,qbar;
assign j=1;
assign k=1;
jk2 jk0(j,k,clk,clr,q[0],qbar[0]);
jk2 jk1(j,k,q[0],clr,q[1],qbar[1]);
jk2 jk3(j,k,q[1],clr,q[2],qbar[2]);
jk2 jk4(j,k,q[2],clr,q[3],qbar[3]);
endmodule
